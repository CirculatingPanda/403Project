//generated per build
//Place a skeleton file here